library ieee;
use ieee.std_logic_1164.all;
use work.eecs361_gates.all;
use work.eecs361.all;

entity control_unit is
  port (
       -- stuff
         );
end control_unit;

architecture structural of control_unit is

        -- component declarations here
begin

        -- logic here

end architecture structural;