library ieee;
use ieee.std_logic_1164.all;
use work.eecs361_gates.all;
use work.eecs361.all;

entity control_unit is
  port (
       instruction  : in  std_logic_vector(31 downto 26);
       
        );
end control_unit;

architecture structural of control_unit is

        -- component declarations here
begin

        -- logic here

end architecture structural;